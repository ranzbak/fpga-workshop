/*
 * Very simple module driving the LED pin low
 */
module led(output o_led_r);

  // Permanent assignments
	assign o_led_r = 1'b0;

endmodule
